/*====================Ports Declaration====================*/
module IF(
 	output reg [31:0] PCin, //address
	output reg [31:0] Instruct, //data
	output reg [31:0] PCout //data
	);

/*====================Variable Declaration====================*/
reg [31:0] aluout; //data

/*====================Function Code====================*/

endmodule