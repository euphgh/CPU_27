/*====================Ports Declaration====================*/
`include "defines.vh"
module ID(
    //sys
	input  wire clk,rst_n,
    input  wire exe_allowin_in,
    output wire id_allowin_out,
    input  wire if_valid_in,
    output wire id_valid_out,
    //datain
 	input wire [31:0] if_PC_in,if_NNPC_in,if_NPC_in, //datar:
    input wire [31:0] if_Instruct_in, //dataw:
	input wire [31:0] wb_wdata_in, //dataw:
	input wire [3:0]  wb_wen_in, //dataw:
    input wire [4:0]  wb_wnum_in, //dataw:
    input wire [2:0] exe_write_type,mem_write_type,wb_write_type, //control{0:wb,1:mem,2:exe,000:nocheck}
    input wire [4:0] exe_wnum,mem_wnum,wb_wnum,
    input wire [31:0] if_NPC_fast_wire,
    input wire  if_exception_in,
    input wire  [4:0]  if_ExcCode_in,
    input wire  [31:0] if_error_VAddr_in,
    input wire  [31:0] wb_cp0_res_in,
    input wire  wb_ClrStpJmp_in,
    //dataout
	output wire [4:0]  id_sel_wbdata_out, //control:
	output wire [1:0]  id_sel_dm_out, //control:
	output wire [31:0] id_RD2_out, //data:
	output wire [12:0] id_aluop_out,
	output wire [31:0] id_aludata1_out, //data:
	output wire [31:0] id_aludata2_out, //data:
    output wire [2:0]  id_sbhw_con_out, //control:
    output wire [4:0]  id_regnum_out,
    output wire [31:0] id_NNPC_out, 
    output wire [31:0] id_PC_out,
    output wire [3:0]  id_addrexc_con_out, //control:地址例外选择子
    output wire [1:0]  id_lr_con_out, //control:onehot模块选择子
    output wire [4:0]  id_lubhw_con_out,
    output wire [2:0] id_write_type_out,
    output wire [7:0] id_mult_div_op,
    output wire [31:0] id_nextPC_out,
    output wire  id_exception_out,
    output wire  id_bd_out,
    output wire  [4:0]  id_ExcCode_out,
    output wire  [7:0]  id_cp0_addr_out,
    output wire  [31:0]  id_error_VAddr_out,
    output wire  id_eret_out,
    output wire  [1:0] id_mftc0_op_out
	);


/*====================Variable Declaration====================*/

//reg Inputs--------------------------------------------------
wire [4:0]  RR1;
wire [4:0]  RR2;
wire [3:0] reg_we ;
wire [4:0]  WR;    
wire [31:0]  WD;
// reg Output
wire [31:0] RD1,RD2;
//------------------------------------------------------------

// signext Inputs---------------------------------------------       
// wire   [15:0]  imm [decoder]
wire   [2:0]  extend_con; //control:选择:imm的符号扩展-0/imm的0扩展-1/off的左移两位扩展-2

// signext Outputs
wire  [31:0]  extend_res;
//------------------------------------------------------------


// decoder Inputs----------------------------------------------      
// decoder Inputs      
wire  [31:0]  Instruct;

// decoder Outputs
wire  [4:0]  rs;
wire  [4:0]  rt;
wire  [4:0]  rd;
wire  [15:0]  imm;
wire  [25:0]  instr_index; 
wire  [4:0]  sa;
wire  [2:0]  sel_wr_con;   
wire  [1:0]  sel_alud1_con;
wire  [1:0]  sel_alud2_con;
// wire  [2:0]  extend_con;[extend]   
wire  [2:0]  bjpc_con;     
wire  [6:0]  brcal_con;    
wire  [12:0]  aluop;       
wire  [2:0]  sbhw_con;     
wire  [1:0]  sel_dm_con;   
wire  [4:0]  sel_wb_con;   
wire  [3:0]  addrexc_con;
wire  [1:0]  lr_con;
wire  [4:0]  lubhw_con;
wire  [1:0]  bjaddrexc_con;
wire  [1:0]  read_type;
wire  [2:0]  write_type;
wire  [7:0]  mult_div_op;
wire  nop;
wire sys_exc,rsvinst_exc,eret,break_exc;
wire [1:0] mftc0_op;
wire [7:0] cp0_addr;
//------------------------------------------------------------

// brcal Inputs ----------------------------------------------       
//wire  [31:0]  RD1; [reg]     
//wire  [31:0]  RD2; [reg]    
//wire  [5:0]  brcal_con; [decoder]
wire [31:0] NPC;
// brcal Outputs
// wire  brcal_out;
//------------------------------------------------------------

// bjpc Inputs-------------------------------------------------
// wire  [31:0]  RD1; [reg]       
// wire  [31:0]  extend_res; [SE]
// wire  [25:0]  instr_index; [decoder]
// wire  [2:0]  bjpc_con; [decorder]   

// bjpc Outputs
wire  [31:0]  bjpc_out;
//------------------------------------------------------------

// others-----------------------------------------------------
wire [31:0] aludata1_wire,aludata2_wire;
wire allowin;
wire ready;
reg valid_r;

wire [31:0] wb_to_id_wdata_w;
wire [3:0] wb_to_id_wen_w ;
wire [4:0] wb_to_id_wnum_w ;

reg  [31:0] if_to_id_PC_r ;
reg  [31:0] if_to_id_NPC_r;
reg  [31:0] if_to_id_NNPC_r ;
reg  [31:0] if_to_id_Instruct_r;
reg  if_to_id_exception_r;
reg  [4:0]  if_to_id_ExcCode_r;
reg  [31:0]  if_to_id_error_VAddr_r;
// wire [4:0] addrexc_con_wire; //control:地址例外选择子[decoder]
// wire [1:0]  lr_con_wire; //control:onehot模块选择子[decoder]
// wire [4:0] lubhw_con_id_wire;[decoder]
wire [31:0] ID_PC;
assign ID_PC = id_PC_out;
wire [4:0] regnum_id_wire;
//------------------------------------------------------------

/*====================Function Code====================*/
always @(posedge clk ) begin
    if (!rst_n||wb_ClrStpJmp_in)begin
       valid_r <= 1'b0; 
    end
    else if (allowin) begin
        valid_r <= if_valid_in ; 
    end
end
assign allowin = !valid_r || (ready && exe_allowin_in)||wb_ClrStpJmp_in;
assign id_allowin_out = allowin;
assign id_valid_out = valid_r && ready;
assign wb_to_id_wdata_w = wb_wdata_in ;
assign wb_to_id_wen_w = wb_wen_in ;
assign wb_to_id_wnum_w = wb_wnum_in ;

always @(posedge clk) begin
    if (!rst_n||(allowin&&(!if_valid_in))||wb_ClrStpJmp_in) begin
        if_to_id_PC_r <= `ini_if_PC_in;
        if_to_id_NPC_r <= `ini_if_NPC_in;
        if_to_id_NNPC_r <= `ini_if_NNPC_in;
        if_to_id_Instruct_r <= `ini_if_Instruct_in;
        if_to_id_exception_r <= `ini_if_exception_in;
        if_to_id_ExcCode_r <= `ini_if_ExcCode_in;
        if_to_id_error_VAddr_r <= `ini_if_error_VAddr_in;
    end
    else if (allowin && if_valid_in) begin
        if_to_id_PC_r <= if_PC_in;
        if_to_id_NPC_r <= if_NPC_in;
        if_to_id_NNPC_r <= if_NNPC_in;
        if_to_id_Instruct_r <= if_Instruct_in;
        if_to_id_exception_r <= if_exception_in;
        if_to_id_ExcCode_r <= if_ExcCode_in;
        if_to_id_error_VAddr_r <= if_error_VAddr_in;
    end
end
Reg  u_Reg (
    .clk                     ( clk      ),
    .rst_n                   ( rst_n    ),
    .reg_we                  ( reg_we   ),
    .RR1                     ( RR1      ),
    .RR2                     ( RR2      ),
    .WR                      ( WR       ),
    .WD                      ( WD       ),

    .RD1                     ( RD1      ),
    .RD2                     ( RD2      )
);
assign id_RD2_out = RD2;
signext  u_signext (
    .imm 		             ( imm		    ),
    .extend_con              ( extend_con   ),

    .extend_res              ( extend_res   ) 
);
decoder  u_decoder (
    .Instruct                ( Instruct        ),

    .rs                      ( rs              ),
    .rt                      ( rt              ),
    .rd                      ( rd              ),
    .imm                     ( imm             ),
    .instr_index             ( instr_index     ),
    .sa                      ( sa              ),
    .sel_wr_con              ( sel_wr_con      ),
    .sel_alud1_con           ( sel_alud1_con   ),
    .sel_alud2_con           ( sel_alud2_con   ),
    .extend_con              ( extend_con      ),
    .bjpc_con                ( bjpc_con        ),
    .brcal_con               ( brcal_con       ),
    .aluop                   ( aluop           ),
    .sbhw_con                ( sbhw_con        ),
    .sel_dm_con              ( sel_dm_con      ),
    .sel_wb_con              ( sel_wb_con      ),
    .addrexc_con             ( addrexc_con     ),
    .lr_con                  ( lr_con          ),
    .lubhw_con               ( lubhw_con       ),
    .read_type               ( read_type       ),
    .write_type              ( write_type      ),
    .mult_div_op             ( mult_div_op     ),
    .nop                     ( nop             ),
    .break_exc               ( break_exc       ),
    .sys_exc                 ( sys_exc         ),
    .mftc0_op                ( mftc0_op        ),
    .eret                    ( eret            ),
    .cp0_addr                ( cp0_addr        ),
    .rsvinst_exc             ( rsvinst_exc     )
);
assign id_sbhw_con_out = sbhw_con;
assign id_lr_con_out = lr_con;
assign id_sel_dm_out = sel_dm_con;
assign id_addrexc_con_out = addrexc_con;
assign id_lubhw_con_out = lubhw_con;
assign id_sel_wbdata_out = sel_wb_con & {5{(!nop)}};
assign Instruct = if_to_id_Instruct_r; //在本阶段没有问题，因为不会出现IF段暂停但是ID段可以继续运行的现象。
assign id_aluop_out = aluop;
assign id_mult_div_op = mult_div_op;
assign regnum_id_wire = sel_wr_con[0] ? rt:
			sel_wr_con[1] ? rd : 32'd31;
assign id_regnum_out = (regnum_id_wire);  //& {5{(!nop)}}) ;
assign aludata1_wire = sel_alud1_con[0] ? RD1 : {27'b0,sa}; //不支持位移负值
assign id_aludata1_out = aludata1_wire;
assign aludata2_wire = sel_alud2_con[0] ? RD2 : extend_res;
assign id_aludata2_out = aludata2_wire;	
assign RR1 = rs;
assign RR2 = rt;
assign WD = wb_to_id_wdata_w;
assign id_PC_out = if_to_id_PC_r;
assign id_NNPC_out = if_to_id_NNPC_r;
assign reg_we = wb_to_id_wen_w; //& {4{valid_r}};
assign WR = wb_to_id_wnum_w;
assign id_write_type_out = write_type & {3{(!nop)}};
idready  u_idready (
    .exe_write_type          ( exe_write_type   ),
    .mem_write_type          ( mem_write_type   ),
    .wb_write_type           ( wb_write_type    ),
    .exe_wnum                ( exe_wnum         ),
    .mem_wnum                ( mem_wnum         ),
    .wb_wnum                 ( wb_wnum          ),
    .read_type               ( read_type        ),
    .RR1                     ( mftc0_op[0] ? rd : RR1  ),
    .RR2                     ( RR2              ),

    .ready                   ( ready            )
);
bjpc  u_bjpc (
    .NPC                     ( NPC           ),
    .RD1                     ( RD1           ),
    .extend_out              ( extend_res    ),
    .instr_index             ( instr_index   ),
    .bjpc_con                ( bjpc_con      ),

    .bjpc_out                ( bjpc_out      )
);
assign NPC = if_to_id_NPC_r;
brcal  u_brcal (
    .RD1                     ( RD1         ),
    .RD2                     ( RD2         ),
    .brcal_con               ( brcal_con   ),

    .brcal_out               ( brcal_out   ) 
);
assign id_nextPC_out = wb_ClrStpJmp_in ? wb_cp0_res_in: (brcal_out ? bjpc_out : if_NPC_fast_wire);
//需要decoder支持
reg bj_last;//表示上一条指令时bj类指令
always @(posedge clk ) begin
    if (!rst_n) 
        bj_last <= 1'b0;
    else
        bj_last <= |brcal_con;
end
assign id_exception_out = if_to_id_exception_r||sys_exc||rsvinst_exc||break_exc;
assign id_bd_out = bj_last;
wire [4:0] ExcCode_id = ({5{rsvinst_exc}} & `RI)|({5{sys_exc}} & `Sys)|({5{break_exc}} & `RI); 
assign id_ExcCode_out = if_to_id_exception_r ? if_to_id_ExcCode_r : ExcCode_id;
assign id_cp0_addr_out = cp0_addr;
assign id_error_VAddr_out = if_to_id_error_VAddr_r;
assign id_eret_out = eret;
assign id_mftc0_op_out = mftc0_op;
endmodule