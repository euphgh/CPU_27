`include "defines.vh"
/*====================Ports Declaration====================*/
module name (
    
    );
/*====================Variable Declaration====================*/

/*====================Function Code====================*/
endmodule