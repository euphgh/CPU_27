`include "defines.vh"
/*====================Ports Declaration====================*/
module alufoward (
    input wire [31:0] alu_res
    
    );
/*====================Variable Declaration====================*/

/*====================Function Code====================*/
endmodule