/*====================Ports Declaration====================*/
module Instr(
 	);

/*====================Variable Declaration====================*/

/*====================Function Code====================*/

endmodule