/*====================Ports Declaration====================*/
module decoder(
 	input wire [31:0] Instruct, //address:

	output wire [4:0] rs, //data:
	output wire [4:0] rt, //data:
	output wire [4:0] rd, //data:
	output wire [15:0] imm, //data:
	output wire [25:0] instr_index, //data:
	output wire [4:0] sa, //data:

	output wire [2:0] sel_wr_con, //control:
	output wire [1:0] sel_alud1_con, //control
	output wire [1:0] sel_alud2_con, //control:
	output wire [2:0] extend_con, //control:
	output wire [2:0] bjpc_con, //control:
	output wire [6:0] brcal_con, //control:
	output wire [12:0] aluop, //control:
	output wire [2:0] sbhw_con, //control:
	output wire [1:0] sel_dm_con, //control:
	output wire [4:0] sel_wb_con, //control:
	output wire [3:0] addrexc_con, //control:地址例外选择子
    output wire [1:0]  lr_con, //control:onehot模块选择子
    output wire [4:0] lubhw_con, //control:lubhw模块选择子
	//new
	output wire [1:0] read_type,
	output wire [2:0] write_type,
	output wire [7:0] mult_div_op,
	output wire nop,
	output wire [1:0] mftc0_op,
	output wire break_exc,
	output wire sys_exc,
	output wire eret,
	output wire [7:0] cp0_addr,
	output wire rsvinst_exc
	);

/*====================Variable Declaration====================*/
wire [31:0] ins = Instruct; 
/*====================Function Code====================*/
//--------------------Manual Code--------------------
assign rs = ins[25:21] ;
assign rt = ins[20:16] ;
assign rd = ins[15:11] ;
assign imm = ins[15:0] ;
assign instr_index = ins[25:0] ;
assign sa = ins[10:6] ;
assign nop = !(|ins);
assign cp0_addr = {ins[15:11],ins[2:0]};
assign rsvinst_exc = !((ins[31:26]==6'd0)||(ins[31:26]==6'd1)||(ins[31:26]==6'd2)||(ins[31:26]==6'd3)||
(ins[31:26]==6'd4)||(ins[31:26]==6'd5)||(ins[31:26]==6'd6)||(ins[31:26]==6'd7)||
(ins[31:26]==6'd8)||(ins[31:26]==6'd9)||(ins[31:26]==6'd10)||(ins[31:26]==6'd11)||
(ins[31:26]==6'd12)||(ins[31:26]==6'd13)||(ins[31:26]==6'd14)||(ins[31:26]==6'd15)||
(ins[31:26]==6'd16)||(ins[31:26]==6'd32)||(ins[31:26]==6'd33)||(ins[31:26]==6'd34)||
(ins[31:26]==6'd35)||(ins[31:26]==6'd36)||(ins[31:26]==6'd37)||(ins[31:26]==6'd38)||
(ins[31:26]==6'd40)||(ins[31:26]==6'd41)||(ins[31:26]==6'd42)||(ins[31:26]==6'd43)||(ins[31:26]==6'd46));
assign write_type[2] = sel_wb_con[3]||sel_wb_con[0];
assign write_type[0] = mftc0_op[0]||sel_wb_con[4];
//--------------------Python Code--------------------
assign break_exc = (!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[3]&&ins[2]&&ins[0] ;
assign sys_exc = (!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[3]&&ins[2]&&(!ins[0]) ;
assign eret = ins[30]&&ins[3] ;
assign mftc0_op[1] = ins[30]&&ins[23];
assign mftc0_op[0] = ins[30]&&(!ins[25])&&(!ins[23]) ;
assign extend_con[0] = (ins[31]||(!ins[29])||(!ins[28])) && (ins[31]||ins[29]||(!ins[28])) && (ins[31]||ins[29]||ins[28]) ;
assign extend_con[1] = ((!ins[31])&&ins[29]&&ins[28]) ;
assign extend_con[2] = ((!ins[31])&&(!ins[29])) ;
assign bjpc_con[0] = ((!ins[31])&&(!ins[28])&&ins[27]) ;
assign bjpc_con[1] = ((!ins[31])&&ins[28]&&(!ins[27])&&(!ins[26])) || ((!ins[31])&&ins[28]&&(!ins[27])&&ins[26]) || ((!ins[31])&&(!ins[28])&&(!ins[27])&&ins[26])
 || ((!ins[31])&&ins[28]&&ins[27]&&ins[26]) || ((!ins[31])&&ins[28]&&ins[27]&&(!ins[26])) ;
assign brcal_con[0] = ((!ins[31])&&(!ins[29])&&ins[28]&&(!ins[27])&&(!ins[26])) ;
assign brcal_con[1] = ((!ins[31])&&(!ins[29])&&ins[28]&&(!ins[27])&&ins[26]) ;
assign brcal_con[3] = ((!ins[29])&&ins[28]&&ins[27]&&ins[26]) ;
assign brcal_con[4] = ((!ins[31])&&(!ins[29])&&ins[28]&&ins[27]&&(!ins[26])) ;
assign sel_alud2_con[1] = (ins[31]||ins[29]||ins[28]||ins[26]) ;
assign aluop[0] = (ins[28]&&ins[27]&&ins[26]) ;
assign sbhw_con[0] = ((!ins[26])) ;
assign sbhw_con[1] = ((!ins[27])&&ins[26]) ;
assign sbhw_con[2] = (ins[27]) ;
assign sel_dm_con[0] = (ins[31]&&ins[29]&&(!ins[27])&&(!ins[26])) || (ins[31]&&ins[29]&&(!ins[27])&&ins[26]) || (ins[31]&&ins[29]&&ins[27]&&ins[26]) ;
assign sel_dm_con[1] = (ins[31]&&ins[29]&&ins[27]&&(!ins[26])) ;
assign sel_wb_con[1] = (ins[31]&&(!ins[29])&&(!ins[27])&&(!ins[26])) || (ins[31]&&(!ins[29])&&(!ins[27])&&ins[26]) || (ins[31]&&(!ins[29])&&ins[27]&&ins[26]) ;
assign sel_wb_con[2] = (ins[31]&&(!ins[29])&&ins[27]&&(!ins[26])) ;
assign addrexc_con[0] = (ins[31]&&(!ins[29])&&(!ins[27])&&ins[26]) ;
assign addrexc_con[1] = (ins[31]&&(!ins[29])&&ins[27]&&ins[26]) ;
assign addrexc_con[2] = (ins[31]&&ins[29]&&(!ins[27])&&ins[26]) ;
assign addrexc_con[3] = (ins[31]&&ins[29]&&ins[27]&&ins[26]) ;
assign lr_con[0] = ((!ins[28])) ;
assign lr_con[1] = (ins[28]) ;
assign lubhw_con[0] = ((!ins[28])&&(!ins[26])) ;
assign lubhw_con[1] = (ins[28]&&(!ins[26])) ;
assign lubhw_con[2] = ((!ins[28])&&(!ins[27])&&ins[26]) ;
assign lubhw_con[3] = (ins[28]&&ins[26]) ;
assign lubhw_con[4] = (ins[27]) ;
assign write_type[1] = (ins[31]&&(!ins[29])) ;
assign bjpc_con[2] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1])) ;
assign brcal_con[2] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[16]) ;
assign brcal_con[5] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&(!ins[16])) ;
assign aluop[10] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&(!ins[3])&&(!ins[2])&&ins[1]) ;
assign aluop[7] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[2]&&ins[1]&&ins[0]) ;
assign aluop[3] = ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[4])&&(!ins[3])&&(!ins[1])) ;
assign aluop[2] = ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[4])&&ins[1]&&(!ins[0])) ;
assign aluop[1] = ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[4])&&ins[1]&&ins[0]) ;
assign sel_wb_con[4] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[0])) ;
assign brcal_con[6] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[2])&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[2])&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[2]&&(!ins[1]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[2]&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[2])&&ins[1])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[2]&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[2]&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[2])&&(!ins[1]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[2])&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[2]&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[2]&&ins[1])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[2])&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[2])&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&ins[2]&&(!ins[1]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&ins[2]&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&(!ins[3])&&(!ins[2])&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&(!ins[3])&&(!ins[2])&&ins[1])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&(!ins[3])&&ins[2]&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&(!ins[3])&&ins[2]&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&ins[3]&&(!ins[2])&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&ins[3]&&ins[2]&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&ins[3]&&ins[2]&&ins[1])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&(!ins[3])&&(!ins[2])&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&(!ins[3])&&(!ins[2])&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&(!ins[3])&&ins[2]&&(!ins[1]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&(!ins[3])&&ins[2]&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&ins[3]&&(!ins[2])&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&ins[3]&&(!ins[2])&&ins[1])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&ins[3]&&ins[2]&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&ins[3]&&ins[2]&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1])) ;
assign sel_wr_con[2] = ((!ins[31])&&(!ins[29])&&ins[26]&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[29])&&ins[26]&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[29])&&ins[26]&&ins[3]&&(!ins[1]))
 || ((!ins[31])&&(!ins[29])&&ins[26]&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[29])&&(!ins[26])&&ins[3]&&(!ins[1])) ;
assign aluop[11] = (ins[31]||ins[29]||ins[28]||ins[27]||(!ins[5])||ins[2]||(!ins[1])) && (ins[31]||(!ins[29])||ins[28]||(!ins[27])||ins[5]||ins[2]||ins[1]) && (ins[31]||(!ins[29])||ins[28]||(!ins[27])||ins[5]||ins[2]||(!ins[1]))
 && (ins[31]||(!ins[29])||ins[28]||(!ins[27])||ins[5]||(!ins[2])||ins[1]) && (ins[31]||(!ins[29])||ins[28]||(!ins[27])||ins[5]||(!ins[2])||(!ins[1])) && (ins[31]||(!ins[29])||ins[28]||(!ins[27])||(!ins[5])||ins[2]||ins[1])
 && (ins[31]||(!ins[29])||ins[28]||(!ins[27])||(!ins[5])||ins[2]||(!ins[1])) && (ins[31]||(!ins[29])||ins[28]||(!ins[27])||(!ins[5])||(!ins[2])||ins[1]) && (ins[31]||(!ins[29])||ins[28]||(!ins[27])||(!ins[5])||(!ins[2])||(!ins[1]))
 && (ins[31]||ins[29]||ins[28]||ins[27]||(!ins[5])||(!ins[2])||ins[1]) && (ins[31]||ins[29]||ins[28]||ins[27]||(!ins[5])||(!ins[2])||(!ins[1])) && (ins[31]||(!ins[29])||(!ins[28])||ins[27]||ins[5]||ins[2]||ins[1])
 && (ins[31]||(!ins[29])||(!ins[28])||ins[27]||ins[5]||ins[2]||(!ins[1])) && (ins[31]||(!ins[29])||(!ins[28])||ins[27]||ins[5]||(!ins[2])||ins[1]) && (ins[31]||(!ins[29])||(!ins[28])||ins[27]||ins[5]||(!ins[2])||(!ins[1]))
 && (ins[31]||(!ins[29])||(!ins[28])||ins[27]||(!ins[5])||ins[2]||ins[1]) && (ins[31]||(!ins[29])||(!ins[28])||ins[27]||(!ins[5])||ins[2]||(!ins[1])) && (ins[31]||(!ins[29])||(!ins[28])||ins[27]||(!ins[5])||(!ins[2])||ins[1])
 && (ins[31]||(!ins[29])||(!ins[28])||ins[27]||(!ins[5])||(!ins[2])||(!ins[1])) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||ins[5]||ins[2]||ins[1]) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||ins[5]||ins[2]||(!ins[1]))
 && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||ins[5]||(!ins[2])||ins[1]) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||ins[5]||(!ins[2])||(!ins[1])) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[5])||ins[2]||ins[1])
 && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[5])||ins[2]||(!ins[1])) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[5])||(!ins[2])||ins[1]) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[5])||(!ins[2])||(!ins[1]))
 && (ins[31]||ins[29]||ins[28]||ins[27]||ins[5]||ins[2]||ins[1]) && (ins[31]||ins[29]||ins[28]||ins[27]||ins[5]||ins[2]||(!ins[1])) && (ins[31]||ins[29]||ins[28]||ins[27]||ins[5]||(!ins[2])||ins[1])
 && (ins[31]||ins[29]||ins[28]||ins[27]||ins[5]||(!ins[2])||(!ins[1])) ;
 assign aluop[9] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[2])&&(!ins[1])&&ins[0])
 || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[5])&&ins[2]&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[5])&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[5])&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[5])&&ins[2]&&ins[1]&&ins[0])
 || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[5]&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[5]&&(!ins[2])&&(!ins[1])&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[5]&&(!ins[2])&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[5]&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[2]&&(!ins[1])&&ins[0])
 || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[2]&&ins[1]&&ins[0]) ;
assign aluop[8] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[2])&&(!ins[1])&&ins[0])
 || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&ins[2]&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&ins[2]&&ins[1]&&ins[0]) ;
assign aluop[6] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[5])&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[5])&&(!ins[2])&&(!ins[1])&&ins[0])
 || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[5])&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[5])&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[5])&&ins[2]&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[5])&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[5])&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[5])&&ins[2]&&ins[1]&&ins[0])
 || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[5]&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[5]&&(!ins[2])&&(!ins[1])&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[5]&&(!ins[2])&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[5]&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[5]&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[5]&&ins[2]&&(!ins[1])&&ins[0])
 || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[5]&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[5]&&ins[2]&&ins[1]&&ins[0]) ;
assign aluop[5] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[3]&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[3])&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[3])&&ins[0])
 || ((!ins[31])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[3]&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[3]&&ins[0]) ;
assign aluop[4] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[3]&&ins[0]) || ((!ins[31])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[3])&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[3])&&ins[0])
 || ((!ins[31])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&ins[3]&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&ins[3]&&ins[0]) ;
assign sel_wb_con[0] = ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&(!ins[4])&&(!ins[3])&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&(!ins[4])&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&(!ins[4])&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&(!ins[4])&&ins[3]&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[4]&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[4]&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[4]&&ins[3]&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[4]&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&ins[3]&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&(!ins[3])&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[4])&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[4])&&(!ins[3])&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[4])&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[4])&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&ins[4]&&(!ins[3])&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&ins[4]&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&ins[4]&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&(!ins[27])&&ins[26]&&ins[4]&&ins[3]&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&ins[26]&&(!ins[4])&&(!ins[3])&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&ins[26]&&(!ins[4])&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&ins[26]&&(!ins[4])&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&ins[26]&&(!ins[4])&&ins[3]&&ins[1])
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&ins[26]&&ins[4]&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&ins[26]&&ins[4]&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&ins[26]&&ins[4]&&ins[3]&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&ins[26]&&ins[4]&&ins[3]&&ins[1]) ;
assign sel_wb_con[3] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&(!ins[2])&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&(!ins[2])&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&ins[2]&&(!ins[1])&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&ins[2]&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&(!ins[2])&&ins[1]&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&ins[2]&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&ins[2]&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&(!ins[2])&&(!ins[1])&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&ins[2]&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&ins[2]&&ins[1]&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&(!ins[2])&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&(!ins[2])&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&ins[2]&&(!ins[1])&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&ins[2]&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&(!ins[3])&&(!ins[2])&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&(!ins[3])&&(!ins[2])&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&(!ins[3])&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&(!ins[3])&&(!ins[2])&&ins[1]&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&(!ins[3])&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&(!ins[3])&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&(!ins[3])&&ins[2]&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&(!ins[3])&&ins[2]&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1])&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&ins[3]&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&ins[3]&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&ins[3]&&ins[2]&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&ins[3]&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&ins[3]&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&(!ins[4])&&ins[3]&&ins[2]&&ins[1]&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&(!ins[3])&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&(!ins[3])&&(!ins[2])&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&(!ins[3])&&(!ins[2])&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&(!ins[3])&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&(!ins[3])&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&(!ins[3])&&ins[2]&&(!ins[1])&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&(!ins[3])&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&(!ins[3])&&ins[2]&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&ins[3]&&(!ins[2])&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&ins[3]&&(!ins[2])&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&ins[3]&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&ins[3]&&(!ins[2])&&ins[1]&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&ins[3]&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&ins[3]&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&ins[3]&&ins[2]&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[20])&&ins[4]&&ins[3]&&ins[2]&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&(!ins[2])&&(!ins[1])&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&ins[2]&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&(!ins[3])&&ins[2]&&ins[1]&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&(!ins[2])&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&ins[2]&&(!ins[1])&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&(!ins[4])&&ins[3]&&ins[2]&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&(!ins[2])&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&(!ins[2])&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&(!ins[2])&&ins[1]&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&ins[2]&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&ins[2]&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&(!ins[3])&&ins[2]&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&(!ins[2])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&(!ins[2])&&(!ins[1])&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&(!ins[2])&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&(!ins[2])&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&ins[2]&&(!ins[1])&&(!ins[0]))
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&ins[2]&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&ins[2]&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[29])&&(!ins[28])&&ins[27]&&ins[26]&&ins[20]&&ins[4]&&ins[3]&&ins[2]&&ins[1]&&ins[0])
 || ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[20])&&(!ins[4])&&ins[3]&&(!ins[2])&&(!ins[1])&&ins[0]) ;
 assign aluop[12] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&(!ins[3])&&(!ins[2])&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[3])&&(!ins[2])&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[3])&&(!ins[2])&&ins[0])
 || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[3])&&ins[2]&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[3])&&ins[2]&&ins[0]) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&ins[3]&&(!ins[2])&&(!ins[0]))
 || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&ins[3]&&(!ins[2])&&ins[0]) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&ins[3]&&ins[2]&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&ins[3]&&ins[2]&&ins[0])
 || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&(!ins[3])&&(!ins[2])&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&(!ins[3])&&(!ins[2])&&ins[0]) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&(!ins[3])&&ins[2]&&(!ins[0]))
 || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&(!ins[3])&&ins[2]&&ins[0]) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[3]&&(!ins[2])&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[3]&&(!ins[2])&&ins[0])
 || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[3]&&ins[2]&&(!ins[0])) || ((!ins[31])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[5]&&ins[3]&&ins[2]&&ins[0]) ;
assign read_type[0] = (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||ins[3]||ins[2]||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||ins[3]||ins[2]||(!ins[0])) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||ins[3]||(!ins[2])||ins[0])
 && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||ins[3]||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||(!ins[3])||ins[2]||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||(!ins[3])||ins[2]||(!ins[0]))
 && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||(!ins[3])||(!ins[2])||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||(!ins[3])||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||ins[3]||ins[2]||ins[0])
 && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||ins[3]||ins[2]||(!ins[0])) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||ins[3]||(!ins[2])||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||ins[3]||(!ins[2])||(!ins[0]))
 && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||(!ins[3])||ins[2]||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||(!ins[3])||ins[2]||(!ins[0])) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||(!ins[3])||(!ins[2])||ins[0])
 && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||(!ins[3])||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||ins[3]||ins[2]||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||ins[3]||ins[2]||(!ins[0]))
 && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||ins[3]||(!ins[2])||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||ins[3]||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||(!ins[3])||ins[2]||ins[0])
 && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||(!ins[3])||ins[2]||(!ins[0])) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||(!ins[3])||(!ins[2])||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||(!ins[3])||(!ins[2])||(!ins[0]))
 && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||ins[3]||ins[2]||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||ins[3]||ins[2]||(!ins[0])) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||ins[3]||(!ins[2])||ins[0])
 && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||ins[3]||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||(!ins[3])||ins[2]||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||(!ins[3])||ins[2]||(!ins[0]))
 && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||(!ins[3])||(!ins[2])||ins[0]) && (ins[31]||ins[30]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||(!ins[3])||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||ins[4]||ins[3]||ins[2]||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||ins[4]||ins[3]||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||ins[4]||ins[3]||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||ins[4]||ins[3]||ins[2]||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||ins[4]||ins[3]||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||ins[4]||ins[3]||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||ins[4]||(!ins[3])||ins[2]||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||ins[4]||(!ins[3])||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||ins[4]||(!ins[3])||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||ins[4]||(!ins[3])||(!ins[2])||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||(!ins[4])||ins[3]||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||(!ins[4])||ins[3]||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||(!ins[4])||ins[3]||(!ins[2])||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||(!ins[4])||ins[3]||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||(!ins[4])||(!ins[3])||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||(!ins[4])||(!ins[3])||ins[2]||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||(!ins[4])||(!ins[3])||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||ins[5]||(!ins[4])||(!ins[3])||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||ins[4]||ins[3]||ins[2]||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||ins[4]||ins[3]||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||ins[4]||ins[3]||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||ins[4]||ins[3]||(!ins[2])||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||ins[4]||(!ins[3])||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||ins[4]||(!ins[3])||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||ins[4]||(!ins[3])||(!ins[2])||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||ins[4]||(!ins[3])||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||(!ins[4])||ins[3]||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||(!ins[4])||ins[3]||ins[2]||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||(!ins[4])||ins[3]||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||(!ins[4])||ins[3]||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||(!ins[4])||(!ins[3])||ins[2]||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||(!ins[4])||(!ins[3])||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||(!ins[4])||(!ins[3])||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||ins[26]||(!ins[5])||(!ins[4])||(!ins[3])||(!ins[2])||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||ins[4]||ins[3]||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||ins[4]||ins[3]||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||ins[4]||ins[3]||(!ins[2])||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||ins[4]||ins[3]||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||ins[4]||(!ins[3])||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||ins[4]||(!ins[3])||ins[2]||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||ins[4]||(!ins[3])||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||ins[4]||(!ins[3])||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||ins[3]||ins[2]||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||ins[3]||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||ins[3]||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||ins[3]||(!ins[2])||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||(!ins[3])||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||(!ins[3])||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||(!ins[3])||(!ins[2])||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||(!ins[3])||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||ins[3]||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||ins[3]||ins[2]||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||ins[3]||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||ins[3]||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||(!ins[3])||ins[2]||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||(!ins[3])||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||(!ins[3])||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||(!ins[3])||(!ins[2])||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||ins[3]||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||ins[3]||ins[2]||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||ins[3]||(!ins[2])||ins[0])
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||ins[3]||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||(!ins[3])||ins[2]||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||(!ins[3])||ins[2]||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||(!ins[3])||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||(!ins[3])||(!ins[2])||(!ins[0])) && (ins[31]||ins[30]||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||ins[4]||(!ins[3])||(!ins[2])||(!ins[0]))
 && (ins[31]||ins[30]||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||ins[4]||(!ins[3])||(!ins[2])||ins[0]) && (ins[31]||ins[30]||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||(!ins[4])||ins[3]||ins[2]||ins[0]) && (ins[31]||(!ins[30])||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||ins[4]||ins[3]||ins[2]||ins[0])
 && (ins[31]||(!ins[30])||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||ins[4]||ins[3]||ins[2]||(!ins[0])) && (ins[31]||(!ins[30])||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||ins[4]||ins[3]||(!ins[2])||ins[0]) && (ins[31]||(!ins[30])||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||ins[4]||ins[3]||(!ins[2])||(!ins[0]))
 && (ins[31]||(!ins[30])||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||(!ins[4])||(!ins[3])||ins[2]||ins[0]) ;
assign sel_wr_con[0] = (ins[31]||ins[30]||ins[29]) ;
assign sel_wr_con[1] = ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])&&ins[0]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]&&(!ins[0]))
 || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]&&ins[0]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1]&&(!ins[0])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1]&&ins[0])
 || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1])&&(!ins[0])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1]&&(!ins[0])) ;
assign sel_alud1_con[1] = ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[5])&&(!ins[4])&&(!ins[3])&&(!ins[2])) ;
assign sel_alud2_con[0] = ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1])
 || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1])) ;
assign sel_alud1_con[0] = (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||ins[3]||ins[2]) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||ins[3]||(!ins[2])) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||(!ins[3])||ins[2])
 && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||ins[4]||(!ins[3])||(!ins[2])) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||ins[3]||ins[2]) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||ins[3]||(!ins[2]))
 && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||(!ins[3])||ins[2]) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||ins[5]||(!ins[4])||(!ins[3])||(!ins[2])) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||ins[3]||ins[2])
 && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||ins[3]||(!ins[2])) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||(!ins[3])||ins[2]) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||ins[4]||(!ins[3])||(!ins[2]))
 && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||ins[3]||ins[2]) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||ins[3]||(!ins[2])) && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||(!ins[3])||ins[2])
 && (ins[31]||(!ins[29])||(!ins[28])||(!ins[27])||(!ins[26])||(!ins[5])||(!ins[4])||(!ins[3])||(!ins[2])) && (ins[31]||ins[29]||ins[28]||ins[27]||ins[26]||ins[5]||ins[4]||ins[3]||ins[2]) ;
assign read_type[1] = ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1])
 || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1])
 || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[4])&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[4])&&(!ins[3])&&ins[1])
 || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[4])&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&ins[26]&&(!ins[4])&&ins[3]&&ins[1]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&ins[26]&&ins[4]&&(!ins[3])&&(!ins[1]))
 || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&ins[26]&&ins[4]&&(!ins[3])&&ins[1]) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&ins[26]&&ins[4]&&ins[3]&&(!ins[1])) || ((!ins[31])&&(!ins[30])&&(!ins[29])&&ins[28]&&(!ins[27])&&ins[26]&&ins[4]&&ins[3]&&ins[1])
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[1]))
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1])
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&(!ins[4])&&(!ins[3])&&(!ins[1]))
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&(!ins[4])&&(!ins[3])&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&(!ins[4])&&ins[3]&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&(!ins[4])&&ins[3]&&ins[1])
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[4]&&(!ins[3])&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[4]&&(!ins[3])&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[4]&&ins[3]&&(!ins[1]))
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&(!ins[27])&&ins[26]&&ins[4]&&ins[3]&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&(!ins[3])&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&(!ins[3])&&ins[1])
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&ins[3]&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&(!ins[4])&&ins[3]&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&(!ins[3])&&(!ins[1]))
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&(!ins[3])&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&ins[3]&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&ins[26]&&ins[4]&&ins[3]&&ins[1])
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[1]))
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1])
 || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&(!ins[28])&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1]))
 || (ins[31]&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&(!ins[4])&&ins[3]&&ins[1])
 || (ins[31]&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1])) || (ins[31]&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1]) || (ins[31]&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1]))
 || (ins[31]&&(!ins[30])&&ins[29]&&ins[28]&&ins[27]&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]) || ((!ins[31])&&ins[30]&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&(!ins[1])) || ((!ins[31])&&ins[30]&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&(!ins[4])&&(!ins[3])&&ins[1]) ;
assign mult_div_op[0] = ((!ins[31])&&(!ins[30])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1])&&(!ins[0])) ;
assign mult_div_op[1] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&(!ins[1])&&ins[0]) ;
assign mult_div_op[2] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]&&(!ins[0])) ;
assign mult_div_op[3] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&ins[3]&&ins[1]&&ins[0]) ;
assign mult_div_op[4] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1])&&(!ins[0])) ;
assign mult_div_op[5] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1]&&(!ins[0])) ;
assign mult_div_op[6] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&(!ins[1])&&ins[0]) ;
assign mult_div_op[7] = ((!ins[31])&&(!ins[29])&&(!ins[28])&&(!ins[27])&&(!ins[26])&&ins[4]&&(!ins[3])&&ins[1]&&ins[0]) ;
endmodule